magic
tech scmos
timestamp 1742847693
<< metal1 >>
rect 0 9052 4 9056
rect 740 8980 744 8984
rect -312 8968 -269 8972
rect -312 8692 -308 8968
rect -148 8960 -144 8962
rect -108 8916 52 8920
rect -4 8768 0 8772
rect -312 8688 -271 8692
rect -312 8404 -308 8688
rect -148 8680 -144 8682
rect -110 8636 52 8640
rect -4 8488 0 8492
rect -312 8400 -265 8404
rect -312 8124 -308 8400
rect -144 8396 -140 8398
rect -104 8352 52 8356
rect -4 8204 0 8208
rect -312 8120 -269 8124
rect -312 7848 -308 8120
rect -144 8112 -140 8114
rect -108 8068 52 8072
rect 0 7928 4 7932
rect -312 7844 -275 7848
rect -312 7572 -308 7844
rect -152 7835 -148 7837
rect -117 7791 52 7795
rect -4 7644 0 7648
rect -312 7568 -277 7572
rect -312 7272 -308 7568
rect -152 7557 -148 7559
rect -117 7513 52 7517
rect -4 7360 0 7364
rect -312 7268 -273 7272
rect -312 6992 -308 7268
rect -148 7260 -144 7262
rect -112 7216 52 7220
rect -4 7076 0 7080
rect -312 6988 -268 6992
rect -312 6704 -308 6988
rect -144 6979 -140 6981
rect -108 6935 52 6939
rect -4 6796 0 6800
rect -312 6700 -274 6704
rect -312 6420 -308 6700
rect -148 6691 -144 6693
rect -113 6647 52 6651
rect -4 6516 0 6520
rect -312 6416 -275 6420
rect -312 6140 -308 6416
rect -152 6411 -148 6413
rect -114 6367 52 6371
rect -4 6236 0 6240
rect -312 6136 -277 6140
rect -312 5860 -308 6136
rect -156 6130 -152 6132
rect -118 6086 52 6090
rect -4 5952 0 5956
rect -312 5856 -277 5860
rect -152 5856 -148 5858
rect -312 5592 -308 5856
rect -116 5812 52 5816
rect -4 5668 0 5672
rect -312 5588 -280 5592
rect -312 5296 -308 5588
rect -156 5575 -152 5577
rect -119 5531 52 5535
rect -4 5388 0 5392
rect -312 5292 -288 5296
rect -312 5020 -308 5292
rect -164 5282 -160 5284
rect -128 5238 52 5242
rect -4 5108 0 5112
rect -312 5016 -288 5020
rect -312 4752 -308 5016
rect -164 5005 -160 5007
rect -129 4961 52 4965
rect -4 4828 0 4832
rect -312 4748 -288 4752
rect -312 4420 -308 4748
rect -168 4736 -164 4738
rect -131 4692 52 4696
rect 0 4524 4 4528
rect -312 4416 -288 4420
rect -312 4148 -308 4416
rect -164 4406 -160 4408
rect -127 4362 52 4366
rect -4 4240 0 4244
rect -312 4144 -287 4148
rect -312 3880 -308 4144
rect -164 4129 -160 4131
rect -126 4085 52 4089
rect -4 3960 0 3964
rect -312 3876 -285 3880
rect -312 3592 -308 3876
rect -160 3864 -156 3866
rect -124 3820 52 3824
rect -4 3676 0 3680
rect -312 3588 -285 3592
rect -312 3328 -308 3588
rect -160 3576 -156 3578
rect -124 3532 52 3536
rect 0 3400 5 3404
rect -312 3324 -293 3328
rect -312 3020 -308 3324
rect -168 3312 -164 3314
rect -132 3268 52 3272
rect -4 3116 0 3120
rect -312 3016 -297 3020
rect -312 2732 -308 3016
rect -172 3009 -168 3011
rect -136 2965 52 2969
rect -4 2832 0 2836
rect -312 2728 -267 2732
rect -312 2464 -308 2728
rect -144 2717 -140 2719
rect -106 2673 52 2677
rect -4 2548 0 2552
rect -312 2460 -268 2464
rect -312 2188 -308 2460
rect -144 2448 -140 2450
rect -108 2404 52 2408
rect -4 2268 0 2272
rect -312 2184 -265 2188
rect -312 1908 -308 2184
rect -140 2168 -136 2170
rect -104 2124 52 2128
rect -4 1988 0 1992
rect -312 1904 -265 1908
rect -312 1636 -308 1904
rect -140 1896 -136 1898
rect -104 1852 52 1856
rect -4 1708 0 1712
rect -312 1632 -265 1636
rect -312 1376 -308 1632
rect -140 1624 -136 1626
rect -104 1580 52 1584
rect -4 1424 0 1428
rect -312 1372 -264 1376
rect -312 1064 -308 1372
rect -140 1360 -136 1362
rect -104 1316 52 1320
rect -4 1140 0 1144
rect -312 1060 -252 1064
rect -312 796 -308 1060
rect -128 1052 -124 1054
rect -91 1008 52 1012
rect -4 860 0 864
rect -312 792 -246 796
rect -312 504 -308 792
rect -124 785 -120 787
rect -86 741 52 745
rect -4 580 0 584
rect -312 500 -246 504
rect -312 220 -308 500
rect -124 491 -120 493
rect -84 447 52 451
rect -4 300 0 304
rect -312 216 -238 220
rect -312 4 -308 216
rect -116 206 -112 208
rect -78 162 52 166
rect -312 0 264 4
<< metal2 >>
rect -108 9016 32 9020
rect -157 8980 4 8984
rect 696 8872 700 8876
rect -112 8736 32 8740
rect -159 8700 4 8704
rect 700 8592 704 8596
rect -107 8452 36 8456
rect -154 8420 4 8424
rect 700 8312 704 8316
rect -108 8168 32 8172
rect -157 8136 4 8140
rect 700 8028 704 8032
rect -117 7891 34 7895
rect -166 7856 4 7860
rect 700 7748 704 7752
rect -117 7613 36 7617
rect -166 7580 8 7584
rect 4 7576 8 7580
rect 700 7468 704 7472
rect -112 7316 32 7320
rect -161 7292 4 7296
rect 700 7184 704 7188
rect -108 7035 36 7039
rect -157 7008 4 7012
rect 700 6900 704 6904
rect -113 6747 36 6751
rect -162 6728 4 6732
rect 700 6620 704 6624
rect -114 6467 35 6471
rect -163 6448 4 6452
rect 700 6340 704 6344
rect -118 6186 36 6190
rect -167 6168 4 6172
rect 700 6060 704 6064
rect -119 5912 35 5916
rect -165 5884 4 5888
rect 700 5776 704 5780
rect -119 5631 35 5635
rect -168 5600 4 5604
rect 692 5492 696 5496
rect -128 5338 33 5342
rect -177 5320 4 5324
rect 700 5212 704 5216
rect -129 5061 36 5065
rect -178 5044 4 5048
rect 772 4932 776 4936
rect -132 4792 33 4796
rect -180 4760 4 4764
rect 768 4652 772 4656
rect -130 4462 35 4466
rect 4 4448 8 4452
rect -176 4444 8 4448
rect 700 4344 704 4348
rect -129 4185 36 4189
rect 4 4168 8 4172
rect -175 4164 8 4168
rect 700 4064 704 4068
rect -129 3920 36 3924
rect -173 3892 4 3896
rect 700 3784 704 3788
rect -130 3632 35 3636
rect -173 3608 4 3612
rect 700 3500 704 3504
rect -132 3368 33 3372
rect -181 3340 8 3344
rect 4 3332 8 3340
rect 700 3220 704 3224
rect -136 3065 32 3069
rect -185 3044 4 3048
rect 700 2940 704 2944
rect -106 2773 32 2777
rect 4 2752 8 2764
rect -155 2748 8 2752
rect 700 2656 704 2660
rect -108 2504 32 2508
rect -157 2480 4 2484
rect 700 2372 704 2376
rect -104 2224 33 2228
rect -153 2200 4 2204
rect 700 2092 704 2096
rect -104 1952 33 1956
rect -153 1920 4 1924
rect 700 1812 704 1816
rect -104 1680 33 1684
rect -153 1652 8 1656
rect 4 1644 8 1652
rect 700 1532 704 1536
rect -104 1436 32 1440
rect -104 1416 -100 1436
rect -153 1388 8 1392
rect 4 1360 8 1388
rect 700 1248 704 1252
rect -91 1108 33 1112
rect -140 1072 4 1076
rect 692 964 696 968
rect -86 841 36 845
rect -135 812 8 816
rect 4 796 8 812
rect 700 684 704 688
rect -85 547 34 551
rect -134 516 4 520
rect 688 404 692 408
rect -78 262 34 266
rect -127 232 8 236
rect 708 124 712 128
<< m2contact >>
rect -161 8980 -157 8984
rect 4 8980 8 8984
rect -112 8916 -108 8920
rect 52 8916 56 8920
rect -163 8700 -159 8704
rect 4 8700 8 8704
rect -116 8636 -110 8640
rect 52 8636 56 8640
rect -158 8420 -154 8424
rect 4 8420 8 8424
rect -108 8352 -104 8356
rect 52 8352 56 8356
rect -161 8136 -157 8140
rect 4 8136 8 8140
rect -112 8068 -108 8072
rect 52 8068 56 8072
rect -170 7856 -166 7860
rect 4 7856 8 7860
rect -124 7791 -117 7795
rect 52 7791 56 7795
rect -170 7580 -166 7584
rect 4 7572 8 7576
rect -124 7513 -117 7517
rect 52 7513 56 7517
rect -165 7292 -161 7296
rect 4 7292 8 7296
rect -116 7216 -112 7220
rect 52 7216 56 7220
rect -161 7008 -157 7012
rect 4 7008 8 7012
rect -112 6935 -108 6939
rect 52 6935 56 6939
rect -166 6728 -162 6732
rect 4 6728 8 6732
rect -120 6647 -113 6651
rect 52 6647 56 6651
rect -167 6448 -163 6452
rect 4 6448 8 6452
rect -120 6367 -114 6371
rect 52 6367 56 6371
rect -171 6168 -167 6172
rect 4 6168 8 6172
rect -124 6086 -118 6090
rect 52 6086 56 6090
rect -169 5884 -165 5888
rect 4 5884 8 5888
rect -120 5812 -116 5816
rect 52 5812 56 5816
rect -172 5600 -168 5604
rect 4 5600 8 5604
rect -124 5531 -119 5535
rect 52 5531 56 5535
rect -181 5320 -177 5324
rect 4 5320 8 5324
rect -132 5238 -128 5242
rect 52 5238 56 5242
rect -182 5044 -178 5048
rect 4 5044 8 5048
rect -136 4961 -129 4965
rect 52 4961 56 4965
rect -184 4760 -180 4764
rect 4 4760 8 4764
rect -136 4692 -131 4696
rect 52 4692 56 4696
rect 4 4452 8 4456
rect -180 4444 -176 4448
rect -132 4362 -127 4366
rect 52 4362 56 4366
rect 4 4172 8 4176
rect -179 4164 -175 4168
rect -132 4085 -126 4089
rect 52 4085 56 4089
rect -177 3892 -173 3896
rect 4 3892 8 3896
rect -128 3820 -124 3824
rect 52 3820 56 3824
rect -177 3608 -173 3612
rect 4 3608 8 3612
rect -128 3532 -124 3536
rect 52 3532 56 3536
rect -185 3340 -181 3344
rect 4 3328 8 3332
rect -136 3268 -132 3272
rect 52 3268 56 3272
rect -189 3044 -185 3048
rect 4 3044 8 3048
rect -140 2965 -136 2969
rect 52 2965 56 2969
rect 4 2764 8 2768
rect -159 2748 -155 2752
rect -112 2673 -106 2677
rect 52 2673 56 2677
rect -161 2480 -157 2484
rect 4 2480 8 2484
rect -112 2404 -108 2408
rect 52 2404 56 2408
rect -157 2200 -153 2204
rect 4 2200 8 2204
rect -108 2124 -104 2128
rect 52 2124 56 2128
rect -157 1920 -153 1924
rect 4 1920 8 1924
rect -108 1852 -104 1856
rect 52 1852 56 1856
rect -157 1652 -153 1656
rect 4 1640 8 1644
rect -108 1580 -104 1584
rect 52 1580 56 1584
rect -157 1388 -153 1392
rect 4 1356 8 1360
rect -108 1316 -104 1320
rect 52 1316 56 1320
rect -144 1072 -140 1076
rect 4 1072 8 1076
rect -96 1008 -91 1012
rect 52 1008 56 1012
rect -139 812 -135 816
rect 4 792 8 796
rect -92 741 -86 745
rect 52 741 56 745
rect -138 516 -134 520
rect 4 516 8 520
rect -88 447 -84 451
rect 52 447 56 451
rect -131 232 -127 236
rect 8 232 12 236
rect -84 162 -78 166
rect 52 162 56 166
use EXC  EXC_0
timestamp 1742590723
transform 1 0 -207 0 1 154
box -32 0 129 112
use EXC  EXC_1
timestamp 1742590723
transform 1 0 -214 0 1 439
box -32 0 129 112
use EXC  EXC_2
timestamp 1742590723
transform 1 0 -215 0 1 733
box -32 0 129 112
use EXC  EXC_3
timestamp 1742590723
transform 1 0 -220 0 1 1000
box -32 0 129 112
use EXC  EXC_4
timestamp 1742590723
transform 1 0 -233 0 1 1308
box -32 0 129 112
use EXC  EXC_5
timestamp 1742590723
transform 1 0 -233 0 1 1572
box -32 0 129 112
use EXC  EXC_6
timestamp 1742590723
transform 1 0 -233 0 1 1844
box -32 0 129 112
use EXC  EXC_7
timestamp 1742590723
transform 1 0 -233 0 1 2116
box -32 0 129 112
use EXC  EXC_8
timestamp 1742590723
transform 1 0 -237 0 1 2396
box -32 0 129 112
use EXC  EXC_9
timestamp 1742590723
transform 1 0 -235 0 1 2665
box -32 0 129 112
use EXC  EXC_10
timestamp 1742590723
transform 1 0 -265 0 1 2957
box -32 0 129 112
use EXC  EXC_11
timestamp 1742590723
transform 1 0 -261 0 1 3260
box -32 0 129 112
use EXC  EXC_12
timestamp 1742590723
transform 1 0 -253 0 1 3524
box -32 0 129 112
use EXC  EXC_13
timestamp 1742590723
transform 1 0 -253 0 1 3812
box -32 0 129 112
use EXC  EXC_14
timestamp 1742590723
transform 1 0 -255 0 1 4077
box -32 0 129 112
use EXC  EXC_15
timestamp 1742590723
transform 1 0 -256 0 1 4354
box -32 0 129 112
use EXC  EXC_16
timestamp 1742590723
transform 1 0 -260 0 1 4684
box -32 0 129 112
use EXC  EXC_17
timestamp 1742590723
transform 1 0 -258 0 1 4953
box -32 0 129 112
use EXC  EXC_18
timestamp 1742590723
transform 1 0 -257 0 1 5230
box -32 0 129 112
use EXC  EXC_19
timestamp 1742590723
transform 1 0 -248 0 1 5523
box -32 0 129 112
use EXC  EXC_20
timestamp 1742590723
transform 1 0 -245 0 1 5804
box -32 0 129 112
use EXC  EXC_21
timestamp 1742590723
transform 1 0 -247 0 1 6078
box -32 0 129 112
use EXC  EXC_22
timestamp 1742590723
transform 1 0 -243 0 1 6359
box -32 0 129 112
use EXC  EXC_23
timestamp 1742590723
transform 1 0 -242 0 1 6639
box -32 0 129 112
use EXC  EXC_24
timestamp 1742590723
transform 1 0 -237 0 1 6927
box -32 0 129 112
use EXC  EXC_25
timestamp 1742590723
transform 1 0 -241 0 1 7208
box -32 0 129 112
use EXC  EXC_26
timestamp 1742590723
transform 1 0 -246 0 1 7505
box -32 0 129 112
use EXC  EXC_27
timestamp 1742590723
transform 1 0 -246 0 1 7783
box -32 0 129 112
use EXC  EXC_28
timestamp 1742590723
transform 1 0 -237 0 1 8060
box -32 0 129 112
use EXC  EXC_29
timestamp 1742590723
transform 1 0 -234 0 1 8344
box -32 0 129 112
use EXC  EXC_30
timestamp 1742590723
transform 1 0 -239 0 1 8628
box -32 0 129 112
use EXC  EXC_31
timestamp 1742590723
transform 1 0 -237 0 1 8908
box -32 0 129 112
use FullAdder32  FullAdder32_0
timestamp 1742755635
transform 1 0 32 0 1 32
box -32 -32 740 9024
<< end >>
