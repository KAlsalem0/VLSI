magic
tech scmos
timestamp 1742739743
<< metal1 >>
rect -60 4400 32 4404
rect -60 4396 -56 4400
rect 28 4392 32 4400
rect -28 4336 16 4340
rect 132 4332 136 4408
rect 424 4336 592 4340
rect 168 4216 176 4220
rect 24 4168 28 4172
rect -36 4164 28 4168
rect 168 4144 172 4216
rect 168 4140 448 4144
rect -56 4116 32 4120
rect 28 4112 32 4116
rect -28 4056 16 4060
rect 132 4052 136 4128
rect 444 4060 448 4140
rect 424 4056 448 4060
rect 168 3936 176 3940
rect 24 3888 28 3892
rect -36 3884 28 3888
rect 168 3864 172 3936
rect 168 3860 452 3864
rect -56 3836 32 3840
rect 28 3832 32 3836
rect -28 3776 16 3780
rect 132 3772 136 3848
rect 448 3780 452 3860
rect 424 3776 452 3780
rect 168 3656 176 3660
rect 24 3608 28 3612
rect -36 3604 28 3608
rect 168 3584 172 3656
rect 168 3580 440 3584
rect -56 3552 32 3556
rect 28 3548 32 3552
rect -28 3492 16 3496
rect 132 3488 136 3564
rect 436 3496 440 3580
rect 424 3492 440 3496
rect 168 3372 176 3376
rect 24 3324 28 3328
rect -36 3320 28 3324
rect 168 3300 172 3372
rect 168 3296 460 3300
rect -56 3276 32 3280
rect 28 3268 32 3276
rect -28 3212 16 3216
rect 132 3208 136 3284
rect 456 3216 460 3296
rect 424 3212 460 3216
rect 168 3092 176 3096
rect 24 3044 28 3048
rect -36 3040 28 3044
rect 168 3020 172 3092
rect 168 3016 444 3020
rect -56 2992 32 2996
rect 28 2988 32 2992
rect -28 2928 16 2932
rect 132 2928 136 3004
rect 440 2936 444 3016
rect 424 2932 444 2936
rect 168 2812 176 2816
rect 24 2764 28 2768
rect -36 2760 28 2764
rect 168 2740 172 2812
rect 168 2736 452 2740
rect -56 2708 32 2712
rect 28 2704 32 2708
rect -28 2648 16 2652
rect 132 2644 136 2720
rect 448 2652 452 2736
rect 424 2648 452 2652
rect 168 2528 176 2532
rect 24 2480 28 2484
rect -36 2476 28 2480
rect 168 2456 172 2528
rect 168 2452 460 2456
rect -56 2424 32 2428
rect 28 2420 32 2424
rect -28 2364 16 2368
rect 132 2360 136 2436
rect 456 2368 460 2452
rect 424 2364 460 2368
rect 168 2244 176 2248
rect 24 2196 28 2200
rect -36 2192 28 2196
rect 168 2172 172 2244
rect 168 2168 452 2172
rect -56 2144 32 2148
rect 28 2140 32 2144
rect -28 2084 16 2088
rect 132 2080 136 2156
rect 448 2088 452 2168
rect 424 2084 452 2088
rect 168 1964 176 1968
rect 24 1916 28 1920
rect -36 1912 28 1916
rect 168 1892 172 1964
rect 168 1888 448 1892
rect -56 1864 32 1868
rect 28 1860 32 1864
rect -28 1804 16 1808
rect 132 1800 136 1876
rect 444 1808 448 1888
rect 424 1804 448 1808
rect 168 1684 176 1688
rect 24 1636 28 1640
rect -36 1632 28 1636
rect 168 1612 172 1684
rect 168 1608 456 1612
rect -56 1584 32 1588
rect 28 1580 32 1584
rect -28 1524 16 1528
rect 132 1520 136 1596
rect 452 1528 456 1608
rect 424 1524 456 1528
rect 168 1404 176 1408
rect 24 1356 28 1360
rect -36 1352 28 1356
rect 168 1332 172 1404
rect 168 1328 456 1332
rect -56 1300 32 1304
rect 28 1296 32 1300
rect -28 1240 16 1244
rect 132 1236 136 1312
rect 452 1244 456 1328
rect 424 1240 456 1244
rect 168 1120 176 1124
rect 24 1072 28 1076
rect -36 1068 28 1072
rect 168 1048 172 1120
rect 168 1044 444 1048
rect -56 1016 32 1020
rect 28 1012 32 1016
rect -28 956 16 960
rect 132 952 136 1028
rect 440 960 444 1044
rect 424 956 444 960
rect 168 836 176 840
rect 24 788 28 792
rect -36 784 28 788
rect 168 764 172 836
rect 168 760 460 764
rect -56 736 32 740
rect 28 732 32 736
rect -28 676 16 680
rect 132 672 136 748
rect 456 680 460 760
rect 424 676 460 680
rect 168 556 176 560
rect 24 508 28 512
rect -36 504 28 508
rect 168 484 172 556
rect 168 480 444 484
rect -56 456 32 460
rect 28 452 32 456
rect -28 400 16 404
rect 132 392 136 468
rect 440 400 444 480
rect 424 396 444 400
rect 168 276 176 280
rect 24 228 28 232
rect -36 224 28 228
rect 168 204 172 276
rect 168 200 436 204
rect -56 176 32 180
rect 28 172 32 176
rect -28 116 16 120
rect 132 112 136 188
rect 432 120 436 200
rect 423 116 436 120
rect 28 -60 32 -48
rect -36 -64 32 -60
rect 172 -84 176 0
<< metal2 >>
rect -60 4120 -56 4392
rect -60 3840 -56 4116
rect -60 3556 -56 3836
rect -60 3280 -56 3552
rect -60 2996 -56 3276
rect -60 2712 -56 2992
rect -60 2428 -56 2708
rect -60 2148 -56 2424
rect -60 1868 -56 2144
rect -60 1588 -56 1864
rect -60 1304 -56 1584
rect -60 1020 -56 1300
rect -60 740 -56 1016
rect -60 460 -56 736
rect -60 180 -56 456
rect -60 -72 -56 176
rect -40 4168 -36 4396
rect 380 4228 588 4232
rect -40 3888 -36 4164
rect 380 3948 588 3952
rect -40 3608 -36 3884
rect 380 3668 588 3672
rect -40 3324 -36 3604
rect 380 3384 588 3388
rect -40 3044 -36 3320
rect 380 3104 588 3108
rect -40 2764 -36 3040
rect 380 2824 588 2828
rect -40 2480 -36 2760
rect 380 2540 588 2544
rect -40 2196 -36 2476
rect 380 2256 588 2260
rect -40 1916 -36 2192
rect 380 1976 588 1980
rect -40 1636 -36 1912
rect 380 1696 588 1700
rect -40 1356 -36 1632
rect 380 1416 588 1420
rect -40 1072 -36 1352
rect 380 1132 588 1136
rect -40 788 -36 1068
rect 380 848 582 852
rect -40 508 -36 784
rect 380 568 588 572
rect -40 228 -36 504
rect 381 288 508 292
rect -40 -60 -36 224
rect 380 8 504 12
rect -40 -72 -36 -64
<< m2contact >>
rect -60 4392 -56 4396
rect 28 4388 32 4392
rect 24 4172 28 4176
rect -40 4164 -36 4168
rect -60 4116 -56 4120
rect 28 4108 32 4112
rect 24 3892 28 3896
rect -40 3884 -36 3888
rect -60 3836 -56 3840
rect 28 3828 32 3832
rect 24 3612 28 3616
rect -40 3604 -36 3608
rect -60 3552 -56 3556
rect 28 3544 32 3548
rect 24 3328 28 3332
rect -40 3320 -36 3324
rect -60 3276 -56 3280
rect 28 3264 32 3268
rect 24 3048 28 3052
rect -40 3040 -36 3044
rect -60 2992 -56 2996
rect 28 2984 32 2988
rect 24 2768 28 2772
rect -40 2760 -36 2764
rect -60 2708 -56 2712
rect 28 2700 32 2704
rect 24 2484 28 2488
rect -40 2476 -36 2480
rect -60 2424 -56 2428
rect 28 2416 32 2420
rect 24 2200 28 2204
rect -40 2192 -36 2196
rect -60 2144 -56 2148
rect 28 2136 32 2140
rect 24 1920 28 1924
rect -40 1912 -36 1916
rect -60 1864 -56 1868
rect 28 1856 32 1860
rect 24 1640 28 1644
rect -40 1632 -36 1636
rect -60 1584 -56 1588
rect 28 1576 32 1580
rect 24 1360 28 1364
rect -40 1352 -36 1356
rect -60 1300 -56 1304
rect 28 1292 32 1296
rect 24 1076 28 1080
rect -40 1068 -36 1072
rect -60 1016 -56 1020
rect 28 1008 32 1012
rect 24 792 28 796
rect -40 784 -36 788
rect -60 736 -56 740
rect 28 728 32 732
rect 24 512 28 516
rect -40 504 -36 508
rect -60 456 -56 460
rect 28 448 32 452
rect 24 232 28 236
rect -40 224 -36 228
rect -60 176 -56 180
rect 28 168 32 172
rect 28 -48 32 -44
rect -40 -64 -36 -60
use FullAdder  FullAdder_0
timestamp 1742590723
transform 1 0 15 0 1 60
box -12 -128 408 112
use FullAdder  FullAdder_1
timestamp 1742590723
transform 1 0 16 0 1 340
box -12 -128 408 112
use FullAdder  FullAdder_2
timestamp 1742590723
transform 1 0 16 0 1 620
box -12 -128 408 112
use FullAdder  FullAdder_3
timestamp 1742590723
transform 1 0 16 0 1 900
box -12 -128 408 112
use FullAdder  FullAdder_4
timestamp 1742590723
transform 1 0 16 0 1 1184
box -12 -128 408 112
use FullAdder  FullAdder_5
timestamp 1742590723
transform 1 0 16 0 1 1468
box -12 -128 408 112
use FullAdder  FullAdder_6
timestamp 1742590723
transform 1 0 16 0 1 1748
box -12 -128 408 112
use FullAdder  FullAdder_7
timestamp 1742590723
transform 1 0 16 0 1 2028
box -12 -128 408 112
use FullAdder  FullAdder_8
timestamp 1742590723
transform 1 0 16 0 1 2308
box -12 -128 408 112
use FullAdder  FullAdder_9
timestamp 1742590723
transform 1 0 16 0 1 2592
box -12 -128 408 112
use FullAdder  FullAdder_10
timestamp 1742590723
transform 1 0 16 0 1 2876
box -12 -128 408 112
use FullAdder  FullAdder_11
timestamp 1742590723
transform 1 0 16 0 1 3156
box -12 -128 408 112
use FullAdder  FullAdder_12
timestamp 1742590723
transform 1 0 16 0 1 3436
box -12 -128 408 112
use FullAdder  FullAdder_13
timestamp 1742590723
transform 1 0 16 0 1 3720
box -12 -128 408 112
use FullAdder  FullAdder_14
timestamp 1742590723
transform 1 0 16 0 1 4000
box -12 -128 408 112
use FullAdder  FullAdder_15
timestamp 1742590723
transform 1 0 16 0 1 4280
box -12 -128 408 112
<< labels >>
rlabel metal1 174 -82 174 -82 1 c
rlabel metal1 -25 118 -25 118 1 b0
rlabel metal1 -25 402 -25 402 1 b1
rlabel metal1 -26 678 -26 678 1 b2
rlabel metal1 -25 958 -25 958 1 b3
rlabel metal1 -26 1242 -26 1242 1 b4
rlabel metal1 -26 1526 -26 1526 1 b5
rlabel metal1 -25 1806 -25 1806 1 b6
rlabel metal1 -25 2085 -25 2085 1 b7
rlabel metal1 -25 2365 -25 2365 1 b8
rlabel metal1 -26 2650 -26 2650 1 b9
rlabel metal1 -26 2930 -26 2930 1 b10
rlabel metal1 -25 3213 -25 3213 1 b11
rlabel metal1 -26 3494 -26 3494 1 b12
rlabel metal1 -25 4058 -25 4058 1 b14
rlabel metal1 -26 4338 -26 4338 1 b15
rlabel metal2 -37 4390 -37 4390 1 gnd
rlabel metal2 -58 4385 -58 4385 3 vdd
rlabel metal1 590 4338 590 4338 7 cout
rlabel metal2 586 4230 586 4230 1 sum15
rlabel metal2 586 3949 586 3949 1 sum14
rlabel metal2 587 3670 587 3670 7 sum13
rlabel metal2 586 3386 586 3386 1 sum12
rlabel metal2 587 3106 587 3106 7 sum11
rlabel metal2 586 2825 586 2825 1 sum10
rlabel metal2 586 2542 586 2542 1 sum9
rlabel metal2 586 2258 586 2258 1 sum8
rlabel metal2 586 1978 586 1978 1 sum7
rlabel metal2 586 1698 586 1698 1 sum6
rlabel metal2 586 1418 586 1418 1 sum5
rlabel metal2 586 1134 586 1134 1 sum4
rlabel metal2 578 850 578 850 1 sum3
rlabel metal2 586 570 586 570 1 sum2
rlabel metal2 506 290 506 290 1 sum1
rlabel metal2 502 10 502 10 1 sum0
rlabel metal1 134 186 134 186 1 a0
rlabel metal1 134 466 134 466 1 a1
rlabel metal1 134 746 134 746 1 a2
rlabel metal1 134 1025 134 1025 1 a3
rlabel metal1 134 1310 134 1310 1 a4
rlabel metal1 134 1593 134 1593 1 a5
rlabel metal1 134 1874 134 1874 1 a6
rlabel metal1 134 2154 134 2154 1 a7
rlabel metal1 134 2434 134 2434 1 a8
rlabel metal1 134 2718 134 2718 1 a9
rlabel metal1 134 3001 134 3001 1 a10
rlabel metal1 135 3282 135 3282 1 a11
rlabel metal1 134 3562 134 3562 1 a12
rlabel metal1 134 3846 134 3846 1 a13
rlabel metal1 134 4126 134 4126 1 a14
rlabel metal1 134 4406 134 4406 5 a15
rlabel metal1 -26 3778 -26 3778 1 b13
<< end >>
