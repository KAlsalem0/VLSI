magic
tech scmos
timestamp 1743079094
<< metal1 >>
rect -12 9060 -8 9064
rect -12 8988 -8 8992
rect 848 8884 852 8992
rect 1584 8988 1588 8992
rect 684 8880 852 8884
rect -16 8776 -12 8780
rect -12 8708 -8 8712
rect 844 8604 848 8712
rect 688 8600 848 8604
rect -16 8496 -12 8500
rect 576 8496 844 8500
rect -12 8428 -8 8432
rect -16 8212 -12 8216
rect -12 8144 -8 8148
rect -12 7936 -8 7940
rect -12 7864 -8 7868
rect 576 7760 580 8496
rect 848 8324 852 8428
rect 688 8320 852 8324
rect 584 8212 844 8216
rect -16 7652 -12 7656
rect -12 7580 -8 7584
rect 584 7480 588 8212
rect 848 8040 852 8144
rect 688 8036 852 8040
rect 592 7936 848 7940
rect -16 7368 -12 7372
rect -12 7300 -8 7304
rect 592 7196 596 7936
rect 848 7760 852 7864
rect 688 7756 852 7760
rect 600 7652 844 7656
rect -16 7084 -12 7088
rect -12 7016 -8 7020
rect 600 6912 604 7652
rect 848 7480 852 7584
rect 688 7476 852 7480
rect 608 7368 844 7372
rect -16 6804 -12 6808
rect -12 6736 -8 6740
rect 608 6632 612 7368
rect 844 7196 848 7304
rect 688 7192 848 7196
rect 616 7084 844 7088
rect -16 6524 -12 6528
rect -12 6456 -8 6460
rect 616 6352 620 7084
rect 848 6912 852 7016
rect 688 6908 852 6912
rect 624 6804 848 6808
rect -16 6244 -12 6248
rect -12 6176 -8 6180
rect 624 6072 628 6804
rect 848 6632 852 6736
rect 688 6628 852 6632
rect 632 6524 844 6528
rect -16 5960 -12 5964
rect -12 5892 -8 5896
rect 632 5788 636 6524
rect 848 6352 852 6456
rect 688 6348 852 6352
rect 640 6244 848 6248
rect -16 5676 -12 5680
rect -12 5608 -8 5612
rect 640 5504 644 6244
rect 848 6072 852 6176
rect 688 6068 852 6072
rect 648 5960 844 5964
rect -16 5396 -12 5400
rect -12 5328 -8 5332
rect 648 5224 652 5960
rect 848 5788 852 5892
rect 688 5784 852 5788
rect 656 5676 844 5680
rect -16 5116 -12 5120
rect -12 5052 -8 5056
rect 656 4944 660 5676
rect 848 5504 852 5608
rect 680 5500 852 5504
rect 664 5396 848 5400
rect -16 4836 -12 4840
rect -12 4768 -8 4772
rect 664 4664 668 5396
rect 848 5224 852 5328
rect 688 5220 852 5224
rect 740 5116 844 5120
rect -12 4532 -8 4536
rect -12 4460 -8 4464
rect 740 4356 744 5116
rect 848 4944 852 5056
rect 760 4940 852 4944
rect 848 4664 852 4772
rect 756 4660 852 4664
rect 848 4356 852 4460
rect 688 4352 852 4356
rect -16 4248 -12 4252
rect 596 4248 844 4252
rect -12 4180 -8 4184
rect -16 3968 -12 3972
rect -12 3900 -8 3904
rect -16 3684 -12 3688
rect -12 3616 -8 3620
rect 596 3512 600 4248
rect 848 4076 852 4184
rect 688 4072 852 4076
rect 604 3968 844 3972
rect -12 3408 -7 3412
rect -12 3336 -8 3340
rect 604 3232 608 3968
rect 848 3796 852 3900
rect 688 3792 768 3796
rect 772 3792 852 3796
rect 612 3684 848 3688
rect -16 3124 -12 3128
rect -12 3052 -8 3056
rect 612 2952 616 3684
rect 844 3512 848 3620
rect 688 3508 848 3512
rect 620 3408 849 3412
rect -16 2840 -12 2844
rect -12 2772 -8 2776
rect 620 2668 624 3408
rect 844 3232 848 3340
rect 688 3228 848 3232
rect 628 3124 844 3128
rect -16 2556 -12 2560
rect -12 2488 -8 2492
rect 628 2384 632 3124
rect 848 2952 852 3052
rect 688 2948 852 2952
rect 640 2840 844 2844
rect -16 2276 -12 2280
rect -12 2208 -8 2212
rect 640 2104 644 2840
rect 848 2668 852 2776
rect 688 2664 852 2668
rect 652 2556 848 2560
rect -16 1996 -12 2000
rect -12 1928 -8 1932
rect 652 1824 656 2556
rect 848 2384 852 2488
rect 688 2380 852 2384
rect 844 2104 848 2212
rect 688 2100 848 2104
rect 848 1824 852 1932
rect 688 1820 852 1824
rect -16 1716 -12 1720
rect -12 1648 -8 1652
rect 684 1648 692 1652
rect 696 1648 852 1652
rect 684 1544 688 1648
rect -16 1432 -12 1436
rect -12 1364 -8 1368
rect 848 1260 852 1368
rect 688 1256 700 1260
rect 704 1256 852 1260
rect -16 1148 -12 1152
rect -12 1080 -8 1084
rect 848 976 852 1084
rect 680 972 708 976
rect 712 972 852 976
rect -16 868 -12 872
rect -12 800 -8 804
rect 684 800 720 804
rect 724 800 848 804
rect 684 696 688 800
rect -16 588 -12 592
rect -12 524 -4 528
rect 848 416 852 524
rect 676 412 732 416
rect 736 412 852 416
rect -16 308 -8 312
rect -8 240 0 244
rect 852 136 856 244
rect 696 132 756 136
rect 760 132 856 136
rect 252 8 1112 12
<< metal2 >>
rect 20 9068 880 9072
rect 20 9048 24 9068
rect 876 9048 880 9068
rect 896 9044 900 9060
rect 1540 8880 1544 8884
rect 1544 8600 1548 8604
rect 1544 8320 1548 8324
rect 1544 8036 1548 8040
rect 1544 7756 1548 7760
rect 1544 7476 1548 7480
rect 1544 7192 1548 7196
rect 1544 6908 1548 6912
rect 1544 6628 1548 6632
rect 1544 6348 1548 6352
rect 1544 6068 1548 6072
rect 1544 5784 1548 5788
rect 1536 5500 1540 5504
rect 1544 5220 1548 5224
rect 1616 4940 1620 4944
rect 768 4532 848 4536
rect 768 3796 772 4532
rect 856 4464 860 4836
rect 1612 4660 1620 4664
rect 1544 4352 1548 4356
rect 1544 4072 1548 4076
rect 1544 3792 1548 3796
rect 1544 3508 1548 3512
rect 1544 3228 1548 3232
rect 1544 2948 1548 2952
rect 1544 2664 1548 2668
rect 1544 2380 1548 2384
rect 692 2276 844 2280
rect 692 1652 696 2276
rect 1544 2100 1548 2104
rect 700 1996 844 2000
rect 700 1260 704 1996
rect 1544 1820 1548 1824
rect 708 1716 844 1720
rect 708 976 712 1716
rect 1544 1540 1548 1544
rect 720 1432 844 1436
rect 720 804 724 1432
rect 1544 1256 1548 1260
rect 732 1148 844 1152
rect 732 416 736 1148
rect 1536 972 1540 976
rect 756 868 844 872
rect 756 136 760 868
rect 1544 692 1548 696
rect 1532 412 1536 416
rect 1552 132 1556 136
rect 40 44 44 56
rect 896 44 900 56
rect 40 40 900 44
<< m2contact >>
rect 896 9060 900 9064
rect 680 8880 684 8884
rect 896 8776 900 8780
rect 684 8600 688 8604
rect 684 8320 688 8324
rect 576 7756 580 7760
rect 684 8036 688 8040
rect 584 7476 588 7480
rect 684 7756 688 7760
rect 592 7192 596 7196
rect 684 7476 688 7480
rect 600 6908 604 6912
rect 684 7192 688 7196
rect 608 6628 612 6632
rect 684 6908 688 6912
rect 616 6348 620 6352
rect 684 6628 688 6632
rect 624 6068 628 6072
rect 684 6348 688 6352
rect 632 5784 636 5788
rect 684 6068 688 6072
rect 640 5500 644 5504
rect 684 5784 688 5788
rect 648 5220 652 5224
rect 676 5500 680 5504
rect 656 4940 660 4944
rect 684 5220 688 5224
rect 664 4660 668 4664
rect 756 4940 760 4944
rect 856 4836 860 4840
rect 752 4660 756 4664
rect 848 4532 852 4536
rect 856 4460 860 4464
rect 684 4352 688 4356
rect 684 4072 688 4076
rect 596 3508 600 3512
rect 684 3792 688 3796
rect 768 3792 772 3796
rect 604 3228 608 3232
rect 684 3508 688 3512
rect 612 2948 616 2952
rect 684 3228 688 3232
rect 620 2664 624 2668
rect 684 2948 688 2952
rect 628 2380 632 2384
rect 684 2664 688 2668
rect 640 2100 644 2104
rect 684 2380 688 2384
rect 844 2276 848 2280
rect 684 2100 688 2104
rect 844 1996 848 2000
rect 652 1820 656 1824
rect 684 1820 688 1824
rect 844 1716 848 1720
rect 692 1648 696 1652
rect 684 1540 688 1544
rect 844 1432 848 1436
rect 684 1256 688 1260
rect 700 1256 704 1260
rect 844 1148 848 1152
rect 676 972 680 976
rect 708 972 712 976
rect 844 868 848 872
rect 720 800 724 804
rect 684 692 688 696
rect 896 588 900 592
rect 672 412 676 416
rect 732 412 736 416
rect 896 308 900 312
rect 692 132 696 136
rect 756 132 760 136
use FullAdder32  FullAdder32_0
timestamp 1742755635
transform 1 0 20 0 1 40
box -32 -32 740 9024
use FullAdder32  FullAdder32_1
timestamp 1742755635
transform 1 0 876 0 1 40
box -32 -32 740 9024
<< labels >>
rlabel metal1 810 10 810 10 1 c
rlabel metal2 802 42 802 42 1 gnd
rlabel metal2 794 9070 794 9070 5 vdd
rlabel metal1 1586 8990 1586 8990 1 cout
rlabel metal1 -6 242 -6 242 1 b0
rlabel metal1 -10 526 -10 526 1 b1
rlabel metal1 -10 802 -10 802 1 b2
rlabel metal1 -10 1082 -10 1082 1 b3
rlabel metal1 -10 1366 -10 1366 1 b4
rlabel metal1 -10 1650 -10 1650 1 b5
rlabel metal1 -10 1930 -10 1930 1 b6
rlabel metal1 -10 2210 -10 2210 1 b7
rlabel metal1 -10 2490 -10 2490 1 b8
rlabel metal1 -10 2774 -10 2774 1 b9
rlabel metal1 -10 3054 -10 3054 1 b10
rlabel metal1 -10 3338 -10 3338 1 b11
rlabel metal1 -10 3618 -10 3618 1 b12
rlabel metal1 -10 3902 -10 3902 1 b13
rlabel metal1 -10 4182 -10 4182 1 b14
rlabel metal1 -10 4462 -10 4462 1 b15
rlabel metal1 -10 4770 -10 4770 1 b16
rlabel metal1 -10 5054 -10 5054 1 b17
rlabel metal1 -10 5330 -10 5330 1 b18
rlabel metal1 -10 5610 -10 5610 1 b19
rlabel metal1 -10 5894 -10 5894 1 b20
rlabel metal1 -10 6178 -10 6178 1 b21
rlabel metal1 -10 6458 -10 6458 1 b22
rlabel metal1 -10 6738 -10 6738 1 b23
rlabel metal1 -10 7018 -10 7018 1 b24
rlabel metal1 -10 7302 -10 7302 1 b25
rlabel metal1 -10 7582 -10 7582 1 b26
rlabel metal1 -10 7866 -10 7866 1 b27
rlabel metal1 -10 8146 -10 8146 1 b28
rlabel metal1 -10 8430 -10 8430 1 b29
rlabel metal1 -10 8710 -10 8710 1 b30
rlabel metal1 -10 8990 -10 8990 1 b31
rlabel metal1 -14 310 -14 310 3 a0
rlabel metal1 -14 590 -14 590 3 a1
rlabel metal1 -14 870 -14 870 3 a2
rlabel metal1 -14 1150 -14 1150 3 a3
rlabel metal1 -14 1434 -14 1434 3 a4
rlabel metal1 -14 1718 -14 1718 3 a5
rlabel metal1 -14 1998 -14 1998 3 a6
rlabel metal1 -14 2278 -14 2278 3 a7
rlabel metal1 -14 2558 -14 2558 3 a8
rlabel metal1 -14 2842 -14 2842 3 a9
rlabel metal1 -14 3126 -14 3126 3 a10
rlabel metal1 -10 3410 -10 3410 1 a11
rlabel metal1 -14 3686 -14 3686 3 a12
rlabel metal1 -14 3970 -14 3970 3 a13
rlabel metal1 -14 4250 -14 4250 3 a14
rlabel metal1 -10 4534 -10 4534 1 a15
rlabel metal1 -14 4838 -14 4838 3 a16
rlabel metal1 -14 5118 -14 5118 3 a17
rlabel metal1 -14 5398 -14 5398 3 a18
rlabel metal1 -14 5678 -14 5678 3 a19
rlabel metal1 -14 5962 -14 5962 3 a20
rlabel metal1 -14 6246 -14 6246 3 a21
rlabel metal1 -14 6526 -14 6526 3 a22
rlabel metal1 -14 6806 -14 6806 3 a23
rlabel metal1 -14 7086 -14 7086 3 a24
rlabel metal1 -14 7370 -14 7370 3 a25
rlabel metal1 -14 7654 -14 7654 3 a26
rlabel metal1 -10 7938 -10 7938 1 a27
rlabel metal1 -14 8214 -14 8214 3 a28
rlabel metal1 -14 8498 -14 8498 3 a29
rlabel metal1 -14 8778 -14 8778 3 a30
rlabel metal1 -10 9062 -10 9062 1 a31
rlabel metal2 1554 134 1554 134 1 sum0
rlabel metal2 1534 414 1534 414 1 sum1
rlabel metal2 1546 694 1546 694 1 sum2
rlabel metal2 1538 974 1538 974 1 sum3
rlabel metal2 1546 1258 1546 1258 1 sum4
rlabel metal2 1546 1542 1546 1542 1 sum5
rlabel metal2 1546 1822 1546 1822 1 sum6
rlabel metal2 1546 2102 1546 2102 1 sum7
rlabel metal2 1546 2382 1546 2382 1 sum8
rlabel metal2 1546 2666 1546 2666 1 sum9
rlabel metal2 1546 2950 1546 2950 1 sum10
rlabel metal2 1546 3230 1546 3230 1 sum11
rlabel metal2 1546 3510 1546 3510 1 sum12
rlabel metal2 1546 3794 1546 3794 1 sum13
rlabel metal2 1546 4074 1546 4074 1 sum14
rlabel metal2 1546 4354 1546 4354 1 sum15
rlabel metal2 1618 4662 1618 4662 7 sum16
rlabel metal2 1618 4942 1618 4942 7 sum17
rlabel metal2 1546 5222 1546 5222 1 sum18
rlabel metal2 1538 5502 1538 5502 1 sum19
rlabel metal2 1546 5786 1546 5786 1 sum20
rlabel metal2 1546 6070 1546 6070 1 sum21
rlabel metal2 1546 6350 1546 6350 1 sum22
rlabel metal2 1546 6630 1546 6630 1 sum23
rlabel metal2 1546 6910 1546 6910 1 sum24
rlabel metal2 1546 7194 1546 7194 1 sum25
rlabel metal2 1546 7478 1546 7478 1 sum26
rlabel metal2 1546 7758 1546 7758 1 sum27
rlabel metal2 1546 8038 1546 8038 1 sum28
rlabel metal2 1546 8322 1546 8322 1 sum29
rlabel metal2 1546 8602 1546 8602 1 sum30
rlabel metal2 1542 8882 1542 8882 1 sum31
<< end >>
