magic
tech scmos
timestamp 1742762006
<< metal1 >>
rect -28 9020 196 9024
rect -28 8948 32 8952
rect 652 8948 708 8952
rect -32 8736 192 8740
rect -28 8668 32 8672
rect -32 8456 192 8460
rect -28 8388 32 8392
rect -32 8172 192 8176
rect -28 8104 32 8108
rect -28 7896 196 7900
rect -28 7824 32 7828
rect -32 7612 192 7616
rect -28 7540 32 7544
rect -32 7328 192 7332
rect -28 7260 32 7264
rect -32 7044 192 7048
rect -28 6976 32 6980
rect -32 6764 192 6768
rect -28 6696 32 6700
rect -32 6484 192 6488
rect -28 6416 32 6420
rect -32 6204 192 6208
rect -28 6136 32 6140
rect -32 5920 192 5924
rect -28 5852 32 5856
rect -32 5636 192 5640
rect -28 5568 32 5572
rect -32 5356 192 5360
rect -28 5288 32 5292
rect -32 5076 192 5080
rect -28 5012 32 5016
rect -32 4796 192 4800
rect -28 4728 32 4732
rect 232 4524 236 4528
rect 232 4520 540 4524
rect -28 4492 196 4496
rect 536 4424 540 4520
rect -28 4420 32 4424
rect -32 4208 192 4212
rect -28 4140 32 4144
rect -32 3928 192 3932
rect -28 3860 32 3864
rect -32 3644 192 3648
rect -28 3576 32 3580
rect -27 3368 197 3372
rect -28 3296 32 3300
rect -32 3084 192 3088
rect -28 3012 32 3016
rect -32 2800 192 2804
rect -28 2732 32 2736
rect -32 2516 192 2520
rect -28 2448 32 2452
rect -32 2236 192 2240
rect -28 2168 32 2172
rect -32 1956 192 1960
rect -28 1888 32 1892
rect -32 1676 192 1680
rect -28 1608 32 1612
rect -32 1392 192 1396
rect -28 1324 32 1328
rect -32 1108 192 1112
rect -28 1040 32 1044
rect -32 828 192 832
rect -28 760 32 764
rect -32 548 192 552
rect -28 484 32 488
rect -32 268 192 272
rect -24 200 36 204
rect 232 -32 236 0
<< metal2 >>
rect 648 8840 664 8844
rect 648 8560 668 8564
rect 648 8280 668 8284
rect 648 7996 668 8000
rect 648 7716 668 7720
rect 648 7436 668 7440
rect 648 7152 668 7156
rect 648 6868 668 6872
rect 648 6588 668 6592
rect 648 6308 668 6312
rect 648 6028 668 6032
rect 648 5744 668 5748
rect 640 5460 660 5464
rect 648 5180 668 5184
rect 568 4900 740 4904
rect 564 4620 736 4624
rect 0 4480 4 4540
rect 20 4480 24 4540
rect 648 4312 668 4316
rect 648 4032 668 4036
rect 648 3752 668 3756
rect 648 3468 668 3472
rect 648 3188 668 3192
rect 648 2908 668 2912
rect 648 2624 668 2628
rect 648 2340 668 2344
rect 648 2060 668 2064
rect 648 1780 668 1784
rect 648 1500 668 1504
rect 648 1216 668 1220
rect 640 932 660 936
rect 648 652 668 656
rect 568 372 676 376
rect 564 92 676 96
use FullAdder16  FullAdder16_0
timestamp 1742739060
transform 1 0 60 0 1 84
box -60 -84 592 4408
use FullAdder16  FullAdder16_1
timestamp 1742739060
transform 1 0 60 0 1 4612
box -60 -84 592 4408
<< labels >>
rlabel metal1 234 -30 234 -30 1 c
rlabel metal1 -22 202 -22 202 1 b0
rlabel metal1 -26 486 -26 486 1 b1
rlabel metal1 -26 762 -26 762 1 b2
rlabel metal1 -26 1042 -26 1042 1 b3
rlabel metal1 -26 1326 -26 1326 1 b4
rlabel metal1 -26 1610 -26 1610 1 b5
rlabel metal1 -26 1890 -26 1890 1 b6
rlabel metal1 -26 2170 -26 2170 1 b7
rlabel metal1 -26 2450 -26 2450 1 b8
rlabel metal1 -26 2734 -26 2734 1 b9
rlabel metal1 -26 3014 -26 3014 1 b10
rlabel metal1 -26 3298 -26 3298 1 b11
rlabel metal1 -26 3577 -26 3577 1 b12
rlabel metal1 -26 3862 -26 3862 1 b13
rlabel metal1 -26 4143 -26 4143 1 b14
rlabel metal1 -26 4423 -26 4423 1 b15
rlabel metal1 -26 4494 -26 4494 1 a15
rlabel metal1 -29 4210 -29 4210 3 a14
rlabel metal1 -30 3930 -30 3930 3 a13
rlabel metal1 -30 3646 -30 3646 3 a12
rlabel metal1 -26 3370 -26 3370 1 a11
rlabel metal1 -30 3086 -30 3086 3 a10
rlabel metal1 -30 2802 -30 2802 3 a9
rlabel metal1 -30 2518 -30 2518 3 a8
rlabel metal1 -30 2239 -30 2239 3 a7
rlabel metal1 -29 1958 -29 1958 3 a6
rlabel metal1 -30 1678 -30 1678 3 a5
rlabel metal1 -30 1394 -30 1394 3 a4
rlabel metal1 -30 1110 -30 1110 3 a3
rlabel metal1 -30 830 -30 830 3 a2
rlabel metal1 -29 550 -29 550 3 a1
rlabel metal1 -30 271 -30 271 3 a0
rlabel metal2 674 94 674 94 1 sum0
rlabel metal2 666 654 666 654 1 sum2
rlabel metal2 658 934 658 934 1 sum3
rlabel metal2 666 1218 666 1218 1 sum4
rlabel metal2 666 1501 666 1501 1 sum5
rlabel metal2 666 1782 666 1782 1 sum6
rlabel metal2 666 2062 666 2062 1 sum7
rlabel metal2 666 2341 666 2341 1 sum8
rlabel metal2 666 2626 666 2626 1 sum9
rlabel metal2 666 2910 666 2910 1 sum10
rlabel metal2 666 3190 666 3190 1 sum11
rlabel metal2 667 3470 667 3470 1 sum12
rlabel metal2 667 3755 667 3755 1 sum13
rlabel metal2 666 4034 666 4034 1 sum14
rlabel metal2 666 4314 666 4314 1 sum15
rlabel metal2 734 4622 734 4622 1 sum16
rlabel metal2 738 4902 738 4902 7 sum17
rlabel metal2 22 4510 22 4510 1 gnd
rlabel metal2 2 4510 2 4510 1 vdd
rlabel metal2 666 5181 666 5181 1 sum18
rlabel metal2 658 5462 658 5462 1 sum19
rlabel metal2 666 5746 666 5746 1 sum20
rlabel metal2 666 6030 666 6030 1 sum21
rlabel metal2 666 6310 666 6310 1 sum22
rlabel metal2 666 6590 666 6590 1 sum23
rlabel metal2 666 6869 666 6869 1 sum24
rlabel metal2 666 7154 666 7154 1 sum25
rlabel metal2 665 7438 665 7438 1 sum26
rlabel metal2 667 7718 667 7718 1 sum27
rlabel metal2 666 7998 666 7998 1 sum28
rlabel metal2 666 8282 666 8282 1 sum29
rlabel metal2 666 8562 666 8562 1 sum30
rlabel metal2 662 8842 662 8842 1 sum31
rlabel metal1 707 8950 707 8950 1 cout
rlabel metal2 674 374 674 374 1 sum1
rlabel metal1 -26 4730 -26 4730 1 b16
rlabel metal1 -26 5014 -26 5014 1 b17
rlabel metal1 -30 4798 -30 4798 3 a16
rlabel metal1 -30 5078 -30 5078 3 a17
rlabel metal1 -26 5290 -26 5290 1 b18
rlabel metal1 -29 5358 -29 5358 3 a18
rlabel metal1 -25 5570 -25 5570 1 b19
rlabel metal1 -30 5638 -30 5638 3 a19
rlabel metal1 -26 5854 -26 5854 1 b20
rlabel metal1 -30 5922 -30 5922 3 a20
rlabel metal1 -26 6138 -26 6138 1 b21
rlabel metal1 -30 6206 -30 6206 3 a21
rlabel metal1 -25 6418 -25 6418 1 b22
rlabel metal1 -30 6486 -30 6486 3 a22
rlabel metal1 -26 6698 -26 6698 1 b23
rlabel metal1 -30 6766 -30 6766 3 a23
rlabel metal1 -26 6978 -26 6978 1 b24
rlabel metal1 -30 7046 -30 7046 3 a24
rlabel metal1 -26 7262 -26 7262 1 b25
rlabel metal1 -30 7330 -30 7330 3 a25
rlabel metal1 -26 7542 -26 7542 1 b26
rlabel metal1 -29 7614 -29 7614 3 a26
rlabel metal1 -26 7826 -26 7826 1 b27
rlabel metal1 -26 7898 -26 7898 1 a27
rlabel metal1 -26 8106 -26 8106 1 b28
rlabel metal1 -29 8174 -29 8174 3 a28
rlabel metal1 -26 8390 -26 8390 1 b29
rlabel metal1 -30 8458 -30 8458 3 a29
rlabel metal1 -26 8670 -26 8670 1 b30
rlabel metal1 -30 8738 -30 8738 3 a30
rlabel metal1 -25 8950 -25 8950 1 b31
rlabel metal1 -26 9022 -26 9022 5 a31
<< end >>
