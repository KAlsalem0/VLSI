magic
tech scmos
timestamp 1743077343
<< metal1 >>
rect 848 8884 852 8992
rect 684 8880 852 8884
rect 844 8604 848 8712
rect 688 8600 848 8604
rect 576 8496 844 8500
rect 576 7760 580 8496
rect 848 8324 852 8428
rect 688 8320 852 8324
rect 584 8212 844 8216
rect 584 7480 588 8212
rect 848 8040 852 8144
rect 688 8036 852 8040
rect 592 7936 848 7940
rect 592 7196 596 7936
rect 848 7760 852 7864
rect 688 7756 852 7760
rect 600 7652 844 7656
rect 600 6912 604 7652
rect 848 7480 852 7584
rect 688 7476 852 7480
rect 608 7368 844 7372
rect 608 6632 612 7368
rect 844 7196 848 7304
rect 688 7192 848 7196
rect 616 7084 844 7088
rect 616 6352 620 7084
rect 848 6912 852 7016
rect 688 6908 852 6912
rect 624 6804 848 6808
rect 624 6072 628 6804
rect 848 6632 852 6736
rect 688 6628 852 6632
rect 632 6524 844 6528
rect 632 5788 636 6524
rect 848 6352 852 6456
rect 688 6348 852 6352
rect 640 6244 848 6248
rect 640 5504 644 6244
rect 848 6072 852 6176
rect 688 6068 852 6072
rect 648 5960 844 5964
rect 648 5224 652 5960
rect 848 5788 852 5892
rect 688 5784 852 5788
rect 656 5676 844 5680
rect 656 4944 660 5676
rect 848 5504 852 5608
rect 680 5500 852 5504
rect 664 5396 848 5400
rect 664 4664 668 5396
rect 848 5224 852 5328
rect 688 5220 852 5224
rect 740 5116 844 5120
rect 740 4356 744 5116
rect 848 4944 852 5056
rect 760 4940 852 4944
rect 848 4664 852 4772
rect 756 4660 852 4664
rect 848 4356 852 4460
rect 688 4352 852 4356
rect 596 4248 844 4252
rect 596 3512 600 4248
rect 848 4076 852 4184
rect 688 4072 852 4076
rect 604 3968 844 3972
rect 604 3232 608 3968
rect 848 3796 852 3900
rect 688 3792 768 3796
rect 772 3792 852 3796
rect 612 3684 848 3688
rect 612 2952 616 3684
rect 844 3512 848 3620
rect 688 3508 848 3512
rect 620 3408 849 3412
rect 620 2668 624 3408
rect 844 3232 848 3340
rect 688 3228 848 3232
rect 628 3124 844 3128
rect 628 2384 632 3124
rect 848 2952 852 3052
rect 688 2948 852 2952
rect 640 2840 844 2844
rect 640 2104 644 2840
rect 848 2668 852 2776
rect 688 2664 852 2668
rect 652 2556 848 2560
rect 652 1824 656 2556
rect 848 2384 852 2488
rect 688 2380 852 2384
rect 844 2104 848 2212
rect 688 2100 848 2104
rect 848 1824 852 1932
rect 688 1820 852 1824
rect 684 1648 692 1652
rect 696 1648 852 1652
rect 684 1544 688 1648
rect 848 1260 852 1368
rect 688 1256 700 1260
rect 704 1256 852 1260
rect 848 976 852 1084
rect 680 972 708 976
rect 712 972 852 976
rect 684 800 720 804
rect 724 800 848 804
rect 684 696 688 800
rect 848 416 852 524
rect 676 412 732 416
rect 736 412 852 416
rect 852 136 856 244
rect 696 132 756 136
rect 760 132 856 136
rect 252 8 1112 12
<< metal2 >>
rect 20 9068 880 9072
rect 20 9048 24 9068
rect 876 9048 880 9068
rect 896 9044 900 9060
rect 768 4532 848 4536
rect 768 3796 772 4532
rect 856 4464 860 4836
rect 692 2276 844 2280
rect 692 1652 696 2276
rect 700 1996 844 2000
rect 700 1260 704 1996
rect 708 1716 844 1720
rect 708 976 712 1716
rect 720 1432 844 1436
rect 720 804 724 1432
rect 732 1148 844 1152
rect 732 416 736 1148
rect 756 868 844 872
rect 756 136 760 868
rect 40 44 44 56
rect 896 44 900 56
rect 40 40 900 44
<< m2contact >>
rect 896 9060 900 9064
rect 680 8880 684 8884
rect 896 8776 900 8780
rect 684 8600 688 8604
rect 684 8320 688 8324
rect 576 7756 580 7760
rect 684 8036 688 8040
rect 584 7476 588 7480
rect 684 7756 688 7760
rect 592 7192 596 7196
rect 684 7476 688 7480
rect 600 6908 604 6912
rect 684 7192 688 7196
rect 608 6628 612 6632
rect 684 6908 688 6912
rect 616 6348 620 6352
rect 684 6628 688 6632
rect 624 6068 628 6072
rect 684 6348 688 6352
rect 632 5784 636 5788
rect 684 6068 688 6072
rect 640 5500 644 5504
rect 684 5784 688 5788
rect 648 5220 652 5224
rect 676 5500 680 5504
rect 656 4940 660 4944
rect 684 5220 688 5224
rect 664 4660 668 4664
rect 756 4940 760 4944
rect 856 4836 860 4840
rect 752 4660 756 4664
rect 848 4532 852 4536
rect 856 4460 860 4464
rect 684 4352 688 4356
rect 684 4072 688 4076
rect 596 3508 600 3512
rect 684 3792 688 3796
rect 768 3792 772 3796
rect 604 3228 608 3232
rect 684 3508 688 3512
rect 612 2948 616 2952
rect 684 3228 688 3232
rect 620 2664 624 2668
rect 684 2948 688 2952
rect 628 2380 632 2384
rect 684 2664 688 2668
rect 640 2100 644 2104
rect 684 2380 688 2384
rect 844 2276 848 2280
rect 684 2100 688 2104
rect 844 1996 848 2000
rect 652 1820 656 1824
rect 684 1820 688 1824
rect 844 1716 848 1720
rect 692 1648 696 1652
rect 684 1540 688 1544
rect 844 1432 848 1436
rect 684 1256 688 1260
rect 700 1256 704 1260
rect 844 1148 848 1152
rect 676 972 680 976
rect 708 972 712 976
rect 844 868 848 872
rect 720 800 724 804
rect 684 692 688 696
rect 896 588 900 592
rect 672 412 676 416
rect 732 412 736 416
rect 896 308 900 312
rect 692 132 696 136
rect 756 132 760 136
use FullAdder32  FullAdder32_0
timestamp 1742755635
transform 1 0 20 0 1 40
box -32 -32 740 9024
use FullAdder32  FullAdder32_1
timestamp 1742755635
transform 1 0 876 0 1 40
box -32 -32 740 9024
<< end >>
