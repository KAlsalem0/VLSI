magic
tech scmos
timestamp 1742755635
<< metal1 >>
rect -28 9020 196 9024
rect -28 8948 32 8952
rect 652 8948 708 8952
rect -32 8736 192 8740
rect -28 8668 32 8672
rect -32 8456 192 8460
rect -28 8388 32 8392
rect -32 8172 192 8176
rect -28 8104 32 8108
rect -28 7896 196 7900
rect -28 7824 32 7828
rect -32 7612 192 7616
rect -28 7540 32 7544
rect -32 7328 192 7332
rect -28 7260 32 7264
rect -32 7044 192 7048
rect -28 6976 32 6980
rect -32 6764 192 6768
rect -28 6696 32 6700
rect -32 6484 192 6488
rect -28 6416 32 6420
rect -32 6204 192 6208
rect -28 6136 32 6140
rect -32 5920 192 5924
rect -28 5852 32 5856
rect -32 5636 192 5640
rect -28 5568 32 5572
rect -32 5356 192 5360
rect -28 5288 32 5292
rect -32 5076 192 5080
rect -28 5012 32 5016
rect -32 4796 192 4800
rect -28 4728 32 4732
rect 232 4524 236 4528
rect 232 4520 540 4524
rect -28 4492 196 4496
rect 536 4424 540 4520
rect -28 4420 32 4424
rect -32 4208 192 4212
rect -28 4140 32 4144
rect -32 3928 192 3932
rect -28 3860 32 3864
rect -32 3644 192 3648
rect -28 3576 32 3580
rect -27 3368 197 3372
rect -28 3296 32 3300
rect -32 3084 192 3088
rect -28 3012 32 3016
rect -32 2800 192 2804
rect -28 2732 32 2736
rect -32 2516 192 2520
rect -28 2448 32 2452
rect -32 2236 192 2240
rect -28 2168 32 2172
rect -32 1956 192 1960
rect -28 1888 32 1892
rect -32 1676 192 1680
rect -28 1608 32 1612
rect -32 1392 192 1396
rect -28 1324 32 1328
rect -32 1108 192 1112
rect -28 1040 32 1044
rect -32 828 192 832
rect -28 760 32 764
rect -32 548 192 552
rect -28 484 32 488
rect -32 268 192 272
rect -24 200 36 204
rect 232 -32 236 0
<< metal2 >>
rect 648 8840 664 8844
rect 648 8560 668 8564
rect 648 8280 668 8284
rect 648 7996 668 8000
rect 648 7716 668 7720
rect 648 7436 668 7440
rect 648 7152 668 7156
rect 648 6868 668 6872
rect 648 6588 668 6592
rect 648 6308 668 6312
rect 648 6028 668 6032
rect 648 5744 668 5748
rect 640 5460 660 5464
rect 648 5180 668 5184
rect 568 4900 740 4904
rect 564 4620 736 4624
rect 0 4480 4 4540
rect 20 4480 24 4540
rect 648 4312 668 4316
rect 648 4032 668 4036
rect 648 3752 668 3756
rect 648 3468 668 3472
rect 648 3188 668 3192
rect 648 2908 668 2912
rect 648 2624 668 2628
rect 648 2340 668 2344
rect 648 2060 668 2064
rect 648 1780 668 1784
rect 648 1500 668 1504
rect 648 1216 668 1220
rect 640 932 660 936
rect 648 652 668 656
rect 568 372 656 376
rect 564 92 676 96
use FullAdder16  FullAdder16_0
timestamp 1742739060
transform 1 0 60 0 1 84
box -60 -84 592 4408
use FullAdder16  FullAdder16_1
timestamp 1742739060
transform 1 0 60 0 1 4612
box -60 -84 592 4408
<< end >>
